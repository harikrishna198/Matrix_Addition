----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/13/2023 03:53:53 PM
-- Design Name: 
-- Module Name: Array_pac - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package array_pac is
type matrix_type2 is array (0 to 1, 0 to 1) of STD_LOGIC_VECTOR (3 downto 0);
end package;


